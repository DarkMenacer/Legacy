//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "20ucs138.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w13;    //: /sn:0 {0}(885,201)(896,201){1}
supply0 w0;    //: /sn:0 {0}(578,264)(578,202){1}
//: {2}(578,198)(578,124){3}
//: {4}(578,120)(578,37)(562,37){5}
//: {6}(576,122)(561,122){7}
//: {8}(576,200)(563,200){9}
supply0 w18;    //: /sn:0 {0}(1028,-100)(1028,-122){1}
reg w10;    //: /sn:0 {0}(639,-92)(655,-92)(655,-58){1}
reg w1;    //: /sn:0 {0}(582,-24)(592,-24)(592,25){1}
//: {2}(590,27)(562,27){3}
//: {4}(592,29)(592,110){5}
//: {6}(590,112)(561,112){7}
//: {8}(592,114)(592,190)(563,190){9}
reg w11;    //: /sn:0 {0}(396,-107)(466,-107)(466,-93){1}
reg w15;    //: /sn:0 {0}(702,4)(725,4){1}
reg [7:0] w9;    //: /sn:0 {0}(#:1177,-10)(1177,-75)(1046,-75){1}
wire w16;    //: /sn:0 {0}(639,-28)(630,-28)(630,213){1}
wire [7:0] w6;    //: /sn:0 {0}(#:523,43)(523,56){1}
//: {2}(525,58)(#:602,58){3}
//: {4}(521,58)(497,58){5}
wire [7:0] w7;    //: /sn:0 {0}(#:694,261)(694,289){1}
//: {2}(696,291)(861,291)(#:861,256){3}
//: {4}(692,291)(673,291){5}
//: {6}(669,291)(445,291)(445,177){7}
//: {8}(447,175)(524,175)(#:524,185){9}
//: {10}(445,173)(445,99){11}
//: {12}(447,97)(522,97)(522,107){13}
//: {14}(445,95)(445,0)(523,0)(#:523,22){15}
//: {16}(671,293)(671,309){17}
wire w34;    //: /sn:0 {0}(793,-14)(749,-14)(749,-9){1}
wire w4;    //: /sn:0 {0}(815,196)(815,201)(837,201){1}
wire [7:0] w25;    //: /sn:0 {0}(#:679,234)(692,234){1}
//: {2}(694,232)(#:694,217){3}
//: {4}(694,236)(#:694,245){5}
wire w22;    //: /sn:0 {0}(759,20)(759,44)(939,44)(939,248)(866,248){1}
wire w36;    //: /sn:0 {0}(485,117)(415,117)(415,-75)(450,-75){1}
wire w3;    //: /sn:0 {0}(639,-16)(635,-16){1}
wire [12:0] w20;    //: /sn:0 {0}(#:799,-29)(876,-29)(876,-73)(#:1011,-73){1}
wire w37;    //: /sn:0 {0}(487,195)(430,195)(430,-63)(450,-63){1}
wire [7:0] w12;    //: /sn:0 {0}(#:638,218)(661,218)(661,147){1}
//: {2}(661,143)(661,60){3}
//: {4}(663,58)(678,58)(678,120){5}
//: {6}(#:680,122)(693,122){7}
//: {8}(697,122)(715,122)(715,57)(877,57)(877,187){9}
//: {10}(695,120)(695,44){11}
//: {12}(678,124)(678,188){13}
//: {14}(659,58)(#:618,58){15}
//: {16}(659,145)(#:627,145){17}
wire [7:0] w19;    //: /sn:0 {0}(#:522,128)(522,143){1}
//: {2}(524,145)(#:611,145){3}
//: {4}(520,145)(498,145){5}
wire w21;    //: /sn:0 {0}(739,20)(739,253)(699,253){1}
wire [1:0] w24;    //: /sn:0 {0}(#:479,-69)(746,-69)(746,-44)(#:793,-44){1}
wire [7:0] w8;    //: /sn:0 {0}(#:793,-24)(777,-24)(777,88){1}
//: {2}(779,90)(803,90){3}
//: {4}(777,92)(777,139){5}
//: {6}(779,141)(845,141)(845,187){7}
//: {8}(775,141)(710,141)(#:710,188){9}
wire [1:0] w17;    //: /sn:0 {0}(668,-34)(#:793,-34){1}
wire w33;    //: /sn:0 {0}(639,-52)(610,-52)(610,53){1}
wire [7:0] w14;    //: /sn:0 {0}(#:524,206)(524,216){1}
//: {2}(526,218)(#:622,218){3}
//: {4}(522,218)(497,218){5}
wire [7:0] w2;    //: /sn:0 {0}(#:861,216)(861,226){1}
//: {2}(859,228)(834,228){3}
//: {4}(861,230)(861,240){5}
wire w5;    //: /sn:0 {0}(486,32)(403,32)(403,-87)(450,-87){1}
wire w38;    //: /sn:0 {0}(450,-51)(435,-51){1}
wire w26;    //: /sn:0 {0}(639,-40)(619,-40)(619,140){1}
//: enddecls

  //: joint g8 (w12) @(661, 58) /w:[ 4 -1 14 3 ]
  //: SWITCH g4 (w11) @(379,-107) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: comment g44 @(511,111) /sn:0
  //: /line:" 1 "
  //: /end
  //: joint g16 (w0) @(578, 200) /w:[ -1 2 8 1 ]
  //: joint g3 (w8) @(777, 141) /w:[ 6 5 8 -1 ]
  //: comment g47 @(840,192) /sn:0
  //: /line:" 1 "
  //: /end
  //: GROUND g17 (w0) @(578,270) /sn:0 /w:[ 0 ]
  //: LED g26 (w14) @(490,218) /sn:0 /R:1 /w:[ 5 ] /type:1
  //: SWITCH g2 (w10) @(622,-92) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: joint g23 (w0) @(578, 122) /w:[ -1 4 6 3 ]
  //: joint g30 (w25) @(694, 234) /w:[ -1 2 1 4 ]
  _GGMUL8 #(124) g1 (.A(w12), .B(w8), .P(w25));   //: @(694,204) /sn:0 /w:[ 13 9 3 ]
  //: joint g24 (w19) @(522, 145) /w:[ 2 1 4 -1 ]
  //: comment g39 @(514,26) /sn:0
  //: /line:" 0 "
  //: /end
  _GGBUFIF8 #(4, 6) g29 (.Z(w7), .I(w25), .E(w21));   //: @(694,251) /sn:0 /R:3 /w:[ 0 5 1 ]
  _GGDECODER2 #(6, 6) g51 (.I(w34), .E(w15), .Z0(w21), .Z1(w22));   //: @(749,4) /sn:0 /w:[ 1 1 0 0 ] /ss:0 /do:0
  _GGBUFIF8 #(4, 6) g18 (.Z(w12), .I(w6), .E(w33));   //: @(608,58) /sn:0 /w:[ 15 3 1 ]
  //: joint g10 (w12) @(661, 145) /w:[ -1 2 16 1 ]
  _GGBUFIF8 #(4, 6) g25 (.Z(w12), .I(w14), .E(w16));   //: @(628,218) /sn:0 /w:[ 0 3 1 ]
  //: LED g49 (w8) @(810,90) /sn:0 /R:3 /w:[ 3 ] /type:1
  _GGREG8 #(10, 10, 20) g6 (.Q(w6), .D(w7), .EN(w0), .CLR(w1), .CK(w5));   //: @(523,32) /sn:0 /w:[ 0 15 5 3 0 ]
  //: DIP g50 (w9) @(1177,1) /sn:0 /R:2 /w:[ 0 ] /st:2 /dn:1
  _GGROM8x13 #(10, 30) g58 (.A(w9), .D(w20), .OE(w18));   //: @(1028,-74) /sn:0 /R:2 /w:[ 1 1 0 ] /mem:"/home/student/Downloads/test.mem"
  //: LED g35 (w4) @(815,189) /sn:0 /w:[ 0 ] /type:0
  //: joint g9 (w12) @(678, 122) /w:[ 6 5 -1 12 ]
  _GGREG8 #(10, 10, 20) g7 (.Q(w19), .D(w7), .EN(w0), .CLR(w1), .CK(w36));   //: @(522,117) /sn:0 /w:[ 0 13 7 7 0 ]
  //: comment g56 @(781,7) /sn:0
  //: /line:" input register"
  //: /line:"   select"
  //: /end
  //: GROUND g59 (w18) @(1028,-128) /sn:0 /R:2 /w:[ 1 ]
  //: LED g22 (w19) @(491,145) /sn:0 /R:1 /w:[ 5 ] /type:1
  //: comment g31 @(967,22) /sn:0
  //: /line:" Instruction Format"
  //: /line:" LSB -> 1 bit op code (1->add, 0->mul)"
  //: /line:"     -> 8 bit D-switch input"
  //: /line:"     -> 2 bit input register selection"
  //: /line:" MSB -> 2 bit output register selection"
  //: /line:""
  //: /line:" Eg:-  01 00 00000001 1"
  //: /line:"      out in d-switch add"
  //: /end
  //: joint g41 (w2) @(861, 228) /w:[ -1 1 2 4 ]
  //: LED g36 (w7) @(671,316) /sn:0 /R:2 /w:[ 17 ] /type:1
  //: joint g33 (w7) @(694, 291) /w:[ 2 1 4 -1 ]
  _GGDECODER4 #(6, 6) g54 (.I(w24), .E(w11), .Z0(w5), .Z1(w36), .Z2(w37), .Z3(w38));   //: @(466,-69) /sn:0 /R:3 /w:[ 0 1 1 1 1 0 ] /ss:0 /do:0
  //: comment g45 @(514,190) /sn:0
  //: /line:" 2 "
  //: /end
  //: LED g42 (w12) @(695,37) /sn:0 /w:[ 11 ] /type:1
  //: LED g40 (w2) @(827,228) /sn:0 /R:1 /w:[ 3 ] /type:1
  assign {w24, w17, w8, w34} = w20; //: CONCAT g52  @(798,-29) /sn:0 /w:[ 1 1 0 0 0 ] /dr:0 /tp:0 /drp:0
  //: LED g12 (w6) @(490,58) /sn:0 /R:1 /w:[ 5 ] /type:1
  //: SWITCH g34 (w13) @(914,201) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  //: joint g28 (w14) @(524, 218) /w:[ 2 1 4 -1 ]
  //: comment g46 @(697,191) /sn:0
  //: /line:" 0 "
  //: /end
  //: comment g57 @(469,-103) /sn:0
  //: /line:" output register"
  //: /line:"   select"
  //: /end
  //: SWITCH g11 (w1) @(565,-24) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: joint g14 (w7) @(445, 175) /w:[ 8 10 -1 7 ]
  //: SWITCH g5 (w15) @(685,4) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: joint g19 (w1) @(592, 27) /w:[ -1 1 2 4 ]
  //: joint g21 (w6) @(523, 58) /w:[ 2 1 4 -1 ]
  _GGBUFIF8 #(4, 6) g32 (.Z(w7), .I(w2), .E(w22));   //: @(861,246) /sn:0 /R:3 /w:[ 3 5 1 ]
  //: joint g20 (w1) @(592, 112) /w:[ -1 5 6 8 ]
  //: joint g43 (w12) @(695, 122) /w:[ 8 10 7 -1 ]
  //: LED g38 (w25) @(672,234) /sn:0 /R:1 /w:[ 0 ] /type:1
  //: joint g15 (w7) @(445, 97) /w:[ 12 14 -1 11 ]
  _GGADD8 #(68, 70, 62, 64) g0 (.A(w8), .B(w12), .S(w2), .CI(w13), .CO(w4));   //: @(861,203) /sn:0 /w:[ 7 9 0 0 1 ]
  _GGBUFIF8 #(4, 6) g27 (.Z(w12), .I(w19), .E(w26));   //: @(617,145) /sn:0 /w:[ 17 3 1 ]
  //: comment g48 @(741,110) /sn:0
  //: /line:" dip-switch input"
  //: /end
  //: joint g37 (w7) @(671, 291) /w:[ 5 -1 6 16 ]
  //: joint g55 (w8) @(777, 90) /w:[ 2 1 -1 4 ]
  _GGREG8 #(10, 10, 20) g13 (.Q(w14), .D(w7), .EN(w0), .CLR(w1), .CK(w37));   //: @(524,195) /sn:0 /w:[ 0 9 9 9 0 ]
  _GGDECODER4 #(6, 6) g53 (.I(w17), .E(w10), .Z0(w33), .Z1(w26), .Z2(w16), .Z3(w3));   //: @(655,-34) /sn:0 /R:3 /w:[ 0 1 0 0 0 0 ] /ss:0 /do:0

endmodule
//: /netlistEnd

