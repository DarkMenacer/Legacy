//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Proj.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w65;    //: /sn:0 {0}(-296,73)(-296,84)(-304,84)(-304,96)(-297,96){1}
supply0 w7;    //: /sn:0 {0}(-212,104)(-212,101)(-221,101){1}
reg w58;    //: /sn:0 {0}(-270,-83)(-270,-78)(-290,-78){1}
supply1 w50;    //: /sn:0 {0}(-788,-233)(-788,-260)(-812,-260){1}
reg w59;    //: /sn:0 {0}(-473,215)(-463,215){1}
reg w62;    //: /sn:0 {0}(-387,210)(-366,210)(-366,206){1}
supply0 w4;    //: /sn:0 {0}(-452,31)(-436,31)(-436,36){1}
reg w56;    //: /sn:0 {0}(-885,-415)(-882,-415)(-882,-388)(-892,-388){1}
supply0 w3;    //: /sn:0 {0}(-378,222)(-378,220)(-387,220){1}
reg [7:0] w60;    //: /sn:0 {0}(#:-639,-421)(-639,-385){1}
supply0 w42;    //: /sn:0 {0}(-894,-324)(-879,-324)(-879,-378)(-892,-378){1}
reg w63;    //: /sn:0 {0}(-210,66)(-208,66)(-208,91)(-221,91){1}
reg w54;    //: /sn:0 {0}(-390,-69)(-390,-73)(-366,-73){1}
reg w84;    //: /sn:0 {0}(-500,-171)(-486,-171){1}
supply0 w21;    //: /sn:0 {0}(-561,-280)(-561,-286)(-660,-286){1}
supply0 w1;    //: /sn:0 {0}(-878,-248)(-878,-263){1}
supply0 w31;    //: /sn:0 {0}(-290,264)(-290,274)(-327,274)(-327,269){1}
reg w53;    //: /sn:0 {0}(-407,28)(-407,21)(-452,21){1}
reg w52;    //: /sn:0 {0}(-549,27)(-549,26)(-528,26){1}
supply0 w2;    //: /sn:0 {0}(-274,-63)(-274,-68)(-290,-68){1}
reg w41;    //: /sn:0 {0}(-987,-265)(-987,-262){1}
reg w85;    //: /sn:0 {0}(-498,-141)(-494,-141)(-494,-153)(-486,-153){1}
reg w55;    //: /sn:0 {0}(-980,-383)(-968,-383){1}
reg w43;    //: /sn:0 {0}(-756,-291)(-736,-291){1}
reg w51;    //: /sn:0 {0}(-564,-298)(-564,-296)(-660,-296){1}
supply0 w40;    //: /sn:0 {0}(-631,-371)(-606,-371)(-606,-349){1}
wire w13;    //: /sn:0 {0}(-752,-10)(-780,-10)(-780,-71){1}
//: {2}(-778,-73)(-751,-73){3}
//: {4}(-782,-73)(-814,-73){5}
//: {6}(-818,-73)(-905,-73)(-905,-84)(-914,-84){7}
//: {8}(-816,-71)(-816,-78){9}
wire [7:0] w6;    //: /sn:0 {0}(-329,-83)(-329,-92)(#:-387,-92)(-387,-107){1}
wire w16;    //: /sn:0 {0}(-914,76)(-828,76){1}
wire [15:0] w34;    //: /sn:0 {0}(#:-699,-301)(-699,-315)(-801,-315){1}
//: {2}(-803,-317)(-803,-344){3}
//: {4}(-805,-315)(#:-831,-315)(-831,-290)(#:-861,-290){5}
wire w88;    //: /sn:0 {0}(-645,-140)(-645,-79)(-570,-79)(-570,-236)(-543,-236){1}
wire w81;    //: /sn:0 {0}(-486,-315)(-514,-315){1}
//: {2}(-516,-317)(-516,-322){3}
//: {4}(-518,-315)(-536,-315)(-536,-66)(-730,-66){5}
wire w25;    //: /sn:0 {0}(-752,10)(-800,10)(-800,-51){1}
//: {2}(-798,-53)(-751,-53){3}
//: {4}(-802,-53)(-873,-53){5}
//: {6}(-877,-53)(-883,-53)(-883,-20)(-914,-20){7}
//: {8}(-875,-51)(-875,-36){9}
wire w39;    //: /sn:0 {0}(-751,-83)(-888,-83)(-888,-114){1}
//: {2}(-886,-116)(-847,-116){3}
//: {4}(-843,-116)(-768,-116)(-768,-20)(-752,-20){5}
//: {6}(-845,-118)(-845,-120)(-845,-120)(-845,-118){7}
//: {8}(-890,-116)(-914,-116){9}
wire [7:0] val;    //: /sn:0 {0}(#:-379,-30)(-379,-40)(-364,-40)(-364,62)(-301,62)(-301,72)(-403,72){1}
//: {2}(-404,72)(-600,72)(-600,-210){3}
//: {4}(-600,-214)(-600,-249){5}
//: {6}(-602,-212)(-749,-212)(-749,-246){7}
wire [1:0] reg0;    //: /sn:0 {0}(#:-360,-259)(-345,-259){1}
//: {2}(-341,-259)(-327,-259)(#:-327,-395)(-545,-395)(-545,-291){3}
//: {4}(-543,-289)(-503,-289){5}
//: {6}(-499,-289)(#:-486,-289){7}
//: {8}(-501,-291)(-501,-292){9}
//: {10}(-545,-287)(#:-545,-204)(-620,-204)(-620,-223){11}
//: {12}(-620,-227)(#:-620,-249){13}
//: {14}(-622,-225)(-704,-225)(-704,-233){15}
//: {16}(-343,-257)(-343,-270){17}
wire [7:0] w22;    //: /sn:0 {0}(#:-424,-441)(-424,-366){1}
//: {2}(#:-422,-364)(-394,-364)(-394,-373){3}
//: {4}(-424,-362)(-424,-344){5}
wire [7:0] w0;    //: /sn:0 {0}(#:-600,52)(-600,61)(-493,61){1}
//: {2}(-491,59)(#:-491,37){3}
//: {4}(-491,63)(-491,69){5}
wire w36;    //: /sn:0 {0}(-751,-78)(-895,-78)(-895,-98){1}
//: {2}(-893,-100)(-831,-100){3}
//: {4}(-827,-100)(-775,-100)(-775,-15)(-752,-15){5}
//: {6}(-829,-102)(-829,-103){7}
//: {8}(-897,-100)(-914,-100){9}
wire [7:0] w20;    //: /sn:0 {0}(#:-359,-30)(-359,-36)(-331,-36){1}
//: {2}(#:-327,-36)(-262,-36){3}
//: {4}(#:-258,-36)(-238,-36)(-238,-42){5}
//: {6}(-260,-34)(-260,86){7}
//: {8}(-329,-38)(#:-329,-62){9}
wire [7:0] w29;    //: /sn:0 {0}(#:-464,-107)(-464,-72){1}
wire w30;    //: /sn:0 {0}(-752,0)(-791,0)(-791,-61){1}
//: {2}(-789,-63)(-751,-63){3}
//: {4}(-793,-63)(-843,-63){5}
//: {6}(-847,-63)(-896,-63)(-896,-52)(-914,-52){7}
//: {8}(-845,-61)(-845,-56){9}
wire [7:0] w12;    //: /sn:0 {0}(#:-484,-72)(-484,-98)(-757,-98)(-757,-218)(-931,-218)(-931,-286){1}
//: {2}(-929,-288)(-896,-288){3}
//: {4}(-931,-290)(-931,-347){5}
//: {6}(-929,-349)(-855,-349)(#:-855,-403)(-671,-403)(-671,-385){7}
//: {8}(-931,-351)(#:-931,-372){9}
//: {10}(-933,-349)(-967,-349){11}
wire [7:0] w19;    //: /sn:0 {0}(#:-475,-43)(-475,-25){1}
//: {2}(#:-477,-23)(-521,-23)(-521,-34){3}
//: {4}(-475,-21)(#:-475,8)(-491,8)(-491,16){5}
wire w18;    //: /sn:0 {0}(-914,44)(-858,44){1}
//: {2}(-854,44)(-751,44){3}
//: {4}(-856,42)(-856,37){5}
wire [7:0] w23;    //: /sn:0 {0}(#:-310,242)(-267,242){1}
//: {2}(-263,242)(-203,242)(-203,240)(-192,240){3}
//: {6}(-190,238)(-190,-496)(-414,-496)(-414,-470){7}
//: {4}(-190,242)(#:-190,252)(-191,252)(-191,254){5}
//: {8}(-265,240)(-265,168)(-223,168)(-223,145){9}
//: {10}(-223,141)(-223,112)(-260,112)(#:-260,107){11}
//: {12}(#:-225,143)(-261,143)(-261,138){13}
wire [3:0] opc;    //: /sn:0 {0}(#:-523,115)(-535,115){1}
//: {2}(-537,113)(-537,93){3}
//: {4}(-539,115)(-657,115)(-657,-197){5}
//: {6}(-655,-199)(-630,-199)(-630,-234){7}
//: {8}(-630,-238)(#:-630,-249){9}
//: {10}(#:-632,-236)(-670,-236)(-670,-246){11}
//: {12}(-659,-199)(-1012,-199)(-1012,-164)(#:-1003,-164){13}
wire w24;    //: /sn:0 {0}(-752,15)(-805,15)(-805,-46){1}
//: {2}(-803,-48)(-751,-48){3}
//: {4}(-807,-48)(-869,-48)(-869,-13)(-887,-13){5}
//: {6}(-891,-13)(-902,-13)(-902,-4)(-914,-4){7}
//: {8}(-889,-11)(-889,-9){9}
wire [7:0] w32;    //: /sn:0 {0}(-434,-470)(-434,-490)(#:-1037,-490)(-1037,244)(-428,244){1}
//: {2}(-424,244)(-345,244){3}
//: {4}(-426,242)(#:-426,226){5}
//: {6}(-426,246)(-426,259){7}
wire w8;    //: /sn:0 {0}(-751,-88)(-881,-88)(-881,-130){1}
//: {2}(-879,-132)(-867,-132){3}
//: {4}(-863,-132)(-766,-132)(-766,-25)(-752,-25){5}
//: {6}(-865,-130)(-865,-136){7}
//: {8}(-883,-132)(-914,-132){9}
wire w46;    //: /sn:0 {0}(-606,-175)(-606,-159){1}
//: {2}(-604,-157)(-576,-157)(-576,-241)(-543,-241){3}
//: {4}(-606,-155)(-606,-135)(-608,-135)(-608,-117){5}
wire w27;    //: /sn:0 {0}(-339,88)(-317,88)(-317,-425)(-460,-425)(-460,-454)(-447,-454){1}
wire w75;    //: /sn:0 {0}(-616,-175)(-616,-165)(-614,-165)(-614,-161){1}
//: {2}(-616,-159)(-645,-159)(-645,-156){3}
//: {4}(-614,-157)(-614,-135)(-613,-135)(-613,-117){5}
wire [7:0] w44;    //: /sn:0 {0}(#:-369,-1)(-369,25){1}
//: {2}(#:-367,27)(-287,27)(-287,17){3}
//: {4}(-369,29)(-369,60)(-382,60)(-382,69){5}
wire w17;    //: /sn:0 {0}(-914,60)(-841,60){1}
//: {2}(-837,60)(-791,60)(-791,49)(-751,49){3}
//: {4}(-839,58)(-839,53)(-839,53)(-839,52){5}
wire w28;    //: /sn:0 {0}(-914,28)(-873,28){1}
//: {2}(-869,28)(-788,28)(-788,39)(-751,39){3}
//: {4}(-871,26)(-871,18){5}
wire w67;    //: /sn:0 {0}(-752,-5)(-785,-5)(-785,-66){1}
//: {2}(-783,-68)(-751,-68){3}
//: {4}(-787,-68)(-825,-68){5}
//: {6}(-829,-68)(-914,-68){7}
//: {8}(-827,-66)(-827,-62)(-827,-62)(-827,-63){9}
wire [7:0] w45;    //: /sn:0 {0}(#:-655,-356)(-655,-343)(-741,-343)(-741,-466)(-931,-466)(#:-931,-393){1}
wire w49;    //: /sn:0 {0}(-914,-148)(-892,-148){1}
//: {2}(-888,-148)(-761,-148)(-761,-30)(-752,-30){3}
//: {4}(-890,-150)(-890,-153){5}
wire [1:0] w78;    //: /sn:0 {0}(#:-403,67)(-403,-207)(-513,-207)(-513,-222)(-503,-222){1}
//: {2}(-499,-222)(-486,-222){3}
//: {4}(-501,-220)(-501,-217){5}
wire [7:0] w11;    //: /sn:0 {0}(#:-426,162)(-426,184){1}
//: {2}(-428,186)(-455,186){3}
//: {4}(-426,188)(-426,205){5}
wire w47;    //: /sn:0 {0}(-611,-96)(-611,-14)(-392,-14){1}
wire w15;    //: /sn:0 {0}(-862,-47)(-862,-56){1}
//: {2}(-860,-58)(-798,-58){3}
//: {4}(-794,-58)(-751,-58){5}
//: {6}(-796,-56)(-796,5)(-752,5){7}
//: {8}(-864,-58)(-890,-58)(-890,-36)(-914,-36){9}
wire w61;    //: /sn:0 {0}(-914,-164)(-906,-164)(-906,-166){1}
wire [15:0] w5;    //: /sn:0 {0}(#:-615,-255)(-615,-258){1}
//: {2}(-613,-260)(-433,-260){3}
//: {4}(-431,-262)(-431,-290){5}
//: {6}(-431,-258)(#:-431,-245){7}
//: {8}(-617,-260)(-641,-260)(-641,-279){9}
//: {10}(#:-639,-281)(-630,-281)(-630,-305){11}
//: {12}(-643,-281)(-654,-281)(-654,-272)(-699,-272)(#:-699,-280){13}
wire w64;    //: /sn:0 {0}(-751,-43)(-867,-43)(-867,12)(-914,12){1}
wire w26;    //: /sn:0 {0}(-324,141)(-339,141){1}
wire [1:0] mode;    //: /sn:0 {0}(#:-723,-223)(-723,-218)(-613,-218){1}
//: {2}(-611,-220)(-611,-240)(-610,-240)(-610,-249){3}
//: {4}(-611,-216)(#:-611,-181){5}
wire w9;    //: /sn:0 {0}(-731,-8)(-339,-8)(-339,-231)(-348,-231){1}
//: {2}(-350,-233)(-350,-237)(-350,-237)(-350,-238){3}
//: {4}(-352,-231)(-360,-231){5}
wire w79;    //: /sn:0 {0}(-522,-238)(-509,-238){1}
//: {2}(-505,-238)(-486,-238){3}
//: {4}(-507,-240)(-507,-244)(-507,-244)(-507,-245){5}
wire w57;    //: /sn:0 {0}(-730,44)(-683,44)(-683,-51){1}
//: {2}(-681,-53)(-588,-53)(-588,-56)(-497,-56){3}
//: {4}(-683,-55)(-683,-371)(-679,-371){5}
//: enddecls

  _GGROM8x16 #(10, 30) g8 (.A(w12), .D(w34), .OE(w1));   //: @(-878,-289) /sn:0 /w:[ 3 5 1 ] /mem:"/home/pranav/Desktop/Computer_Science/TkGate/rom.mem"
  _GGMUX2x8 #(8, 8) g4 (.I0(val), .I1(w20), .S(w47), .Z(w44));   //: @(-369,-14) /sn:0 /w:[ 0 0 1 0 ] /ss:0 /do:0
  //: joint g116 (opc) @(-537, 115) /w:[ 1 2 4 -1 ]
  //: LED g17 (w16) @(-821,76) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: joint g137 (w5) @(-431, -260) /w:[ -1 4 3 6 ]
  //: joint g92 (w18) @(-856, 44) /w:[ 2 4 1 -1 ]
  //: joint g74 (w39) @(-845, -116) /w:[ 4 6 3 -1 ]
  //: joint g30 (opc) @(-657, -199) /w:[ 6 -1 12 5 ]
  //: joint g130 (reg0) @(-620, -225) /w:[ -1 12 14 11 ]
  _GGROM8x8 #(10, 30) g1 (.A(w32), .D(w23), .OE(w31));   //: @(-327,243) /sn:0 /w:[ 3 0 1 ] /mem:"/home/pranav/Desktop/Computer_Science/TkGate/rom.mem"
  //: LED g77 (w13) @(-816,-85) /sn:0 /w:[ 9 ] /type:0
  _GGREG8 #(10, 10, 20) PC (.Q(w12), .D(w45), .EN(w42), .CLR(w56), .CK(w55));   //: @(-931,-383) /w:[ 9 1 1 1 1 ]
  //: LED g111 (w44) @(-287,10) /sn:0 /w:[ 3 ] /type:1
  //: SWITCH g51 (w58) @(-270,-96) /sn:0 /R:3 /w:[ 0 ] /st:1 /dn:0
  //: joint g70 (w49) @(-890, -148) /w:[ 2 4 1 -1 ]
  ALU g10 (.in1(w0), .in2(w44), .opc(opc), .ALU_out(w11), .LD(w27), .ST(w26));   //: @(-522, 70) /sz:(182, 91) /sn:0 /p:[ Ti0>5 Ti1>5 Li0>0 Bo0<0 Ro0<0 Ro1<1 ]
  assign {w75, w46} = mode; //: CONCAT g25  @(-611,-180) /sn:0 /R:1 /w:[ 0 0 5 ] /dr:0 /tp:0 /drp:0
  //: joint g65 (w15) @(-796, -58) /w:[ 4 -1 3 6 ]
  //: LED g103 (w78) @(-501,-210) /sn:0 /R:2 /w:[ 5 ] /type:1
  //: joint g64 (w30) @(-791, -63) /w:[ 2 -1 4 1 ]
  //: joint g72 (w8) @(-865, -132) /w:[ 4 -1 3 6 ]
  //: SWITCH g49 (w54) @(-390,-55) /sn:0 /R:1 /w:[ 0 ] /st:1 /dn:0
  //: joint g136 (w5) @(-615, -260) /w:[ 2 -1 8 1 ]
  //: joint g6 (w32) @(-426, 244) /w:[ 2 4 1 6 ]
  //: LED g7 (w34) @(-803,-351) /sn:0 /w:[ 3 ] /type:1
  //: LED g124 (w22) @(-394,-380) /sn:0 /w:[ 3 ] /type:1
  //: joint g58 (reg0) @(-545, -289) /w:[ 4 3 -1 10 ]
  //: SWITCH g56 (w63) @(-227,66) /sn:0 /w:[ 0 ] /st:0 /dn:0
  assign w78 = val[1:0]; //: TAP g35 @(-403,70) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:0
  //: joint g98 (w79) @(-507, -238) /w:[ 2 4 1 -1 ]
  //: LED g85 (w25) @(-875,-29) /sn:0 /R:2 /w:[ 9 ] /type:0
  //: joint g67 (w24) @(-805, -48) /w:[ 2 -1 4 1 ]
  //: joint g126 (w34) @(-803, -315) /w:[ 1 2 4 -1 ]
  //: SWITCH g54 (w62) @(-366,193) /sn:0 /R:3 /w:[ 1 ] /st:1 /dn:0
  _GGAND2 #(6) g33 (.I0(w46), .I1(w88), .Z(w79));   //: @(-532,-238) /sn:0 /w:[ 3 1 0 ]
  //: joint g81 (w30) @(-845, -63) /w:[ 5 -1 6 8 ]
  //: SWITCH g52 (w59) @(-490,215) /sn:0 /w:[ 0 ] /st:1 /dn:0
  //: joint g40 (w57) @(-683, -53) /w:[ 2 4 -1 1 ]
  //: LED g132 (mode) @(-723,-230) /sn:0 /w:[ 0 ] /type:1
  //: VDD g12 (w50) @(-799,-233) /sn:0 /R:2 /w:[ 0 ]
  //: joint g108 (w19) @(-475, -23) /w:[ -1 1 2 4 ]
  //: joint g131 (mode) @(-611, -218) /w:[ -1 2 1 4 ]
  //: joint g106 (reg0) @(-343, -259) /w:[ 2 -1 1 16 ]
  //: joint g96 (w81) @(-516, -315) /w:[ 1 2 4 -1 ]
  assign {opc, reg0, mode, val} = w5; //: CONCAT g19  @(-615,-254) /sn:0 /R:1 /w:[ 9 13 3 5 0 ] /dr:0 /tp:0 /drp:0
  //: joint g114 (w0) @(-491, 61) /w:[ -1 2 1 4 ]
  //: LED g117 (w11) @(-462,186) /sn:0 /R:1 /w:[ 3 ] /type:1
  //: joint g125 (w22) @(-424, -364) /w:[ 2 1 -1 4 ]
  //: joint g78 (w13) @(-816, -73) /w:[ 5 -1 6 8 ]
  //: LED g93 (w17) @(-839,45) /sn:0 /w:[ 5 ] /type:0
  //: joint g63 (w67) @(-785, -68) /w:[ 2 -1 4 1 ]
  //: joint g100 (w9) @(-350, -231) /w:[ 1 2 4 -1 ]
  //: LED g105 (reg0) @(-343,-277) /sn:0 /w:[ 17 ] /type:1
  //: LED g113 (w0) @(-600,45) /sn:0 /w:[ 0 ] /type:1
  //: GROUND g38 (w1) @(-878,-242) /sn:0 /w:[ 0 ]
  //: GROUND g43 (w21) @(-561,-274) /sn:0 /w:[ 0 ]
  _GGMUX2x8 #(8, 8) g0 (.I0(w32), .I1(w23), .S(w27), .Z(w22));   //: @(-424,-454) /sn:0 /w:[ 0 7 1 0 ] /ss:0 /do:0
  //: LED g101 (reg0) @(-501,-299) /sn:0 /w:[ 9 ] /type:1
  //: SWITCH g48 (w53) @(-407,42) /sn:0 /R:1 /w:[ 0 ] /st:1 /dn:0
  _GGREG8 #(10, 10, 20) Rz (.Q(w32), .D(w11), .EN(w3), .CLR(w62), .CK(w59));   //: @(-426,215) /w:[ 5 5 1 0 1 ]
  _GGOR3 #(8) g37 (.I0(w28), .I1(w18), .I2(w17), .Z(w57));   //: @(-740,44) /sn:0 /w:[ 3 3 3 0 ]
  //: joint g80 (w67) @(-827, -68) /w:[ 5 -1 6 8 ]
  //: LED g95 (w81) @(-516,-329) /sn:0 /w:[ 3 ] /type:0
  //: LED g120 (w23) @(-261,131) /sn:0 /w:[ 13 ] /type:1
  //: LED g122 (w23) @(-191,261) /sn:0 /R:2 /w:[ 5 ] /type:1
  //: joint g76 (w36) @(-829, -100) /w:[ 4 6 3 -1 ]
  //: LED g75 (w36) @(-829,-110) /sn:0 /w:[ 7 ] /type:0
  //: SWITCH g44 (w43) @(-773,-291) /sn:0 /w:[ 0 ] /st:1 /dn:0
  //: GROUND g47 (w4) @(-436,42) /sn:0 /w:[ 1 ]
  //: joint g16 (w12) @(-931, -349) /w:[ 6 8 10 5 ]
  //: GROUND g3 (w31) @(-290,258) /sn:0 /R:2 /w:[ 0 ]
  //: joint g90 (w28) @(-871, 28) /w:[ 2 4 1 -1 ]
  _GGXOR2 #(8) g26 (.I0(w46), .I1(w75), .Z(w47));   //: @(-611,-106) /sn:0 /R:3 /w:[ 5 5 0 ]
  _GGREG16 #(10, 10, 20) IR (.Q(w5), .D(w34), .EN(w21), .CLR(w51), .CK(w43));   //: @(-699,-291) /w:[ 13 0 1 1 1 ]
  //: LED g109 (w20) @(-238,-49) /sn:0 /w:[ 5 ] /type:1
  //: joint g2 (w23) @(-190, 240) /w:[ -1 6 3 4 ]
  //: joint g128 (opc) @(-630, -236) /w:[ -1 8 10 7 ]
  //: joint g23 (w12) @(-931, -288) /w:[ 2 4 -1 1 ]
  //: LED g91 (w18) @(-856,30) /sn:0 /w:[ 5 ] /type:0
  //: LED g127 (opc) @(-670,-253) /sn:0 /w:[ 11 ] /type:1
  //: joint g86 (w25) @(-875, -53) /w:[ 5 -1 6 8 ]
  _GGMUX2x8 #(8, 8) g39 (.I0(w29), .I1(w12), .S(w57), .Z(w19));   //: @(-474,-56) /sn:0 /w:[ 1 0 3 0 ] /ss:0 /do:1
  dec4to16 g24 (.opc(opc), .o0(w61), .o1(w49), .o2(w8), .o3(w39), .o4(w36), .o5(w13), .o6(w67), .o7(w30), .o8(w15), .o9(w25), .o10(w24), .o11(w64), .o12(w28), .o13(w18), .o14(w17), .o15(w16));   //: @(-1002, -180) /sz:(87, 272) /sn:0 /p:[ Li0>13 Ro0<0 Ro1<0 Ro2<9 Ro3<9 Ro4<9 Ro5<7 Ro6<7 Ro7<7 Ro8<9 Ro9<7 Ro10<7 Ro11<1 Ro12<0 Ro13<0 Ro14<0 Ro15<0 ]
  //: joint g104 (w78) @(-501, -222) /w:[ 2 -1 1 4 ]
  //: joint g60 (w39) @(-888, -116) /w:[ 2 -1 8 1 ]
  //: SWITCH g29 (w85) @(-515,-141) /sn:0 /w:[ 0 ] /st:0 /dn:0
  _GGREG8 #(10, 10, 20) Rm (.Q(w23), .D(w20), .EN(w7), .CLR(w63), .CK(w65));   //: @(-260,96) /w:[ 11 7 1 1 1 ]
  //: joint g110 (w20) @(-260, -36) /w:[ 4 -1 3 6 ]
  //: joint g121 (w23) @(-223, 143) /w:[ -1 10 12 9 ]
  //: LED g82 (w30) @(-845,-49) /sn:0 /R:2 /w:[ 9 ] /type:0
  //: DIP g18 (w60) @(-639,-431) /sn:0 /w:[ 0 ] /st:4 /dn:0
  //: joint g94 (w17) @(-839, 60) /w:[ 2 4 1 -1 ]
  //: LED g119 (w32) @(-426,266) /sn:0 /R:2 /w:[ 7 ] /type:1
  //: LED g107 (w19) @(-521,-41) /sn:0 /w:[ 3 ] /type:1
  //: GROUND g50 (w2) @(-274,-57) /sn:0 /w:[ 0 ]
  //: LED g133 (val) @(-749,-253) /sn:0 /w:[ 7 ] /type:1
  //: LED g73 (w39) @(-845,-125) /sn:0 /w:[ 7 ] /type:0
  //: joint g9 (w20) @(-329, -36) /w:[ 2 8 1 -1 ]
  _GGREG8 #(10, 10, 20) Ra (.Q(w0), .D(w19), .EN(w4), .CLR(w53), .CK(w52));   //: @(-491,26) /w:[ 3 5 0 1 1 ]
  //: LED g68 (w12) @(-974,-349) /sn:0 /R:1 /w:[ 11 ] /type:1
  //: LED g71 (w8) @(-865,-143) /sn:0 /w:[ 7 ] /type:0
  _GGOR10 #(22) g59 (.I0(w49), .I1(w8), .I2(w39), .I3(w36), .I4(w13), .I5(w67), .I6(w30), .I7(w15), .I8(w25), .I9(w24), .Z(w9));   //: @(-741,-8) /sn:0 /w:[ 3 5 5 5 0 0 0 7 0 0 0 ]
  _GGNBUF #(2) g31 (.I(w75), .Z(w88));   //: @(-645,-150) /sn:0 /R:3 /w:[ 3 0 ]
  //: SWITCH g22 (w56) @(-902,-415) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: joint g102 (reg0) @(-501, -289) /w:[ 6 8 5 -1 ]
  //: LED g87 (w24) @(-889,-2) /sn:0 /R:2 /w:[ 9 ] /type:0
  //: joint g83 (w15) @(-862, -58) /w:[ 2 -1 8 1 ]
  //: LED g99 (w9) @(-350,-245) /sn:0 /w:[ 3 ] /type:0
  //: SWITCH g45 (w51) @(-564,-311) /sn:0 /R:3 /w:[ 0 ] /st:1 /dn:0
  //: LED g41 (w61) @(-906,-173) /sn:0 /w:[ 1 ] /type:0
  _GGOR10 #(22) g36 (.I0(w8), .I1(w39), .I2(w36), .I3(w13), .I4(w67), .I5(w30), .I6(w15), .I7(w25), .I8(w24), .I9(w64), .Z(w81));   //: @(-740,-66) /sn:0 /w:[ 0 0 0 3 3 3 5 3 3 0 5 ]
  //: LED g138 (w5) @(-630,-312) /sn:0 /w:[ 11 ] /type:1
  //: LED g69 (w49) @(-890,-160) /sn:0 /w:[ 5 ] /type:0
  //: joint g42 (w8) @(-881, -132) /w:[ 2 -1 8 1 ]
  //: joint g66 (w25) @(-800, -53) /w:[ 2 -1 4 1 ]
  //: SWITCH g57 (w65) @(-296,60) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH g46 (w52) @(-549,41) /sn:0 /R:1 /w:[ 0 ] /st:1 /dn:0
  //: joint g34 (w46) @(-606, -157) /w:[ 2 1 -1 4 ]
  //: SWITCH g28 (w84) @(-517,-171) /sn:0 /w:[ 0 ] /st:1 /dn:0
  //: joint g5 (w23) @(-265, 242) /w:[ 2 8 1 -1 ]
  //: LED g84 (w15) @(-862,-40) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: GROUND g14 (w42) @(-900,-324) /sn:0 /R:3 /w:[ 0 ]
  //: joint g118 (w11) @(-426, 186) /w:[ -1 1 2 4 ]
  //: joint g112 (w44) @(-369, 27) /w:[ 2 1 -1 4 ]
  //: joint g61 (w36) @(-895, -100) /w:[ 2 -1 8 1 ]
  //: SWITCH g21 (w55) @(-997,-383) /sn:0 /w:[ 0 ] /st:1 /dn:0
  //: joint g32 (w75) @(-614, -159) /w:[ -1 1 2 4 ]
  //: LED g115 (opc) @(-537,86) /sn:0 /w:[ 3 ] /type:1
  //: GROUND g20 (w40) @(-606,-343) /sn:0 /w:[ 1 ]
  //: LED g79 (w67) @(-827,-56) /sn:0 /R:2 /w:[ 9 ] /type:0
  //: joint g134 (val) @(-600, -212) /w:[ -1 4 6 3 ]
  //: LED g97 (w79) @(-507,-252) /sn:0 /w:[ 5 ] /type:0
  //: LED g129 (reg0) @(-704,-240) /sn:0 /w:[ 15 ] /type:1
  //: LED g89 (w28) @(-871,11) /sn:0 /w:[ 5 ] /type:0
  _GGADD8 #(68, 70, 62, 64) g15 (.A(w12), .B(w60), .S(w45), .CI(w40), .CO(w57));   //: @(-655,-369) /sn:0 /w:[ 7 1 0 0 5 ]
  Reg_file g27 (.C(w22), .CLR(w85), .CLK(w84), .Rb_s(w78), .en_Rb(w79), .Ra_s(reg0), .en_Ra(w81), .Rc_s(reg0), .en_Rc(w9), .toRb(w6), .toRa(w29));   //: @(-485, -343) /sz:(124, 235) /sn:0 /p:[ Ti0>5 Li0>1 Li1>1 Li2>3 Li3>3 Li4>7 Li5>0 Ri0>0 Ri1>5 Bo0<1 Bo1<0 ]
  //: joint g62 (w13) @(-780, -73) /w:[ 2 -1 4 1 ]
  //: joint g88 (w24) @(-889, -13) /w:[ 5 -1 6 8 ]
  //: GROUND g55 (w7) @(-212,110) /sn:0 /w:[ 0 ]
  //: LED g135 (w5) @(-431,-297) /sn:0 /w:[ 5 ] /type:1
  _GGREG8 #(10, 10, 20) Rb (.Q(w20), .D(w6), .EN(w2), .CLR(w58), .CK(w54));   //: @(-329,-73) /w:[ 9 0 1 1 1 ]
  //: SWITCH g13 (w41) @(-987,-248) /sn:0 /R:1 /w:[ 1 ] /st:0 /dn:0
  //: GROUND g53 (w3) @(-378,228) /sn:0 /w:[ 0 ]
  //: joint g139 (w5) @(-641, -281) /w:[ 10 -1 12 9 ]

endmodule
//: /netlistEnd

//: /netlistBegin ALU
module ALU(in2, opc, LD, ALU_out, ST, in1);
//: interface  /sz:(182, 91) /bd:[ Ti0>in2[7:0](140/182) Ti1>in1[7:0](31/182) Li0>opc[3:0](45/91) Bo0<ALU_out[7:0](96/182) Ro0<ST(71/91) Ro1<LD(18/91) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply0 w4;    //: /sn:0 {0}(315,202)(315,212)(345,212)(345,217){1}
supply0 w3;    //: /sn:0 {0}(314,114)(314,118)(313,118)(313,133){1}
output LD;    //: /sn:0 {0}(531,-4)(531,42)(550,42){1}
input [7:0] in1;    //: {0}(#:111,127)(120,127){1}
//: {2}(124,127)(129,127){3}
//: {4}(133,127)(-62:138,127)(138,74)(#:300,74){5}
//: {6}(131,129)(131,160){7}
//: {8}(133,162)(301,162){9}
//: {10}(131,164)(131,237){11}
//: {12}(133,239)(#:300,239){13}
//: {14}(131,241)(131,315){15}
//: {16}(133,317)(295,317){17}
//: {18}(131,319)(131,383){19}
//: {20}(133,385)(301,385){21}
//: {22}(#:131,387)(131,413){23}
//: {24}(133,415)(303,415){25}
//: {26}(131,417)(131,441)(#:307,441){27}
//: {28}(122,129)(122,467)(324,467){29}
output [7:0] ALU_out;    //: /sn:0 {0}(#:443,88)(649,88){1}
//: {2}(651,86)(651,71)(650,71)(#:650,55){3}
//: {4}(651,90)(651,132)(650,132)(650,174){5}
//: {6}(648,176)(#:427,176){7}
//: {8}(650,178)(650,251){9}
//: {10}(648,253)(#:411,253){11}
//: {12}(650,255)(650,319){13}
//: {14}(648,321)(#:395,321){15}
//: {16}(650,323)(650,339){17}
//: {18}(648,341)(#:369,341){19}
//: {20}(650,343)(650,379){21}
//: {22}(648,381)(#:389,381){23}
//: {24}(650,383)(650,409){25}
//: {26}(648,411)(#:372,411){27}
//: {28}(650,413)(650,436){29}
//: {30}(648,438)(#:360,438){31}
//: {32}(650,440)(650,465)(#:340,465){33}
output ST;    //: /sn:0 {0}(515,-4)(515,58)(552,58){1}
input [3:0] opc;    //: /sn:0 {0}(#:531,-93)(531,-127)(532,-127)(532,-129){1}
input [7:0] in2;    //: /sn:0 {0}(#:303,410)(142,410)(142,382){1}
//: {2}(144,380)(301,380){3}
//: {4}(142,378)(#:142,351){5}
//: {6}(144,349)(#:295,349){7}
//: {8}(142,347)(142,273){9}
//: {10}(144,271)(#:300,271){11}
//: {12}(142,269)(142,196){13}
//: {14}(144,194)(186,194){15}
//: {16}(140,194)(139,194)(139,149){17}
//: {18}(141,147)(180,147)(180,106)(300,106){19}
//: {20}(137,147)(#:112,147){21}
wire w13;    //: /sn:0 {0}(451,-4)(451,368)(381,368)(381,378){1}
wire [7:0] w6;    //: /sn:0 {0}(301,194)(#:202,194){1}
wire w22;    //: /sn:0 {0}(307,-4)(307,11){1}
wire w0;    //: /sn:0 {0}(315,154)(315,150)(349,150)(349,135){1}
wire w20;    //: /sn:0 {0}(339,-4)(339,11){1}
wire [7:0] o1;    //: /sn:0 {0}(#:324,413)(356,413){1}
wire [7:0] o5;    //: /sn:0 {0}(#:329,255)(395,255){1}
wire [7:0] w37;    //: /sn:0 {0}(#:324,343)(353,343){1}
wire w19;    //: /sn:0 {0}(355,-4)(355,11){1}
wire w18;    //: /sn:0 {0}(371,-4)(371,323)(361,323)(361,338){1}
wire w12;    //: /sn:0 {0}(467,-4)(467,400)(364,400)(364,408){1}
wire w23;    //: /sn:0 {0}(291,-4)(291,11){1}
wire [7:0] o0;    //: /sn:0 {0}(#:323,441)(324,441)(324,440)(344,440){1}
wire w21;    //: /sn:0 {0}(323,-4)(323,11){1}
wire [7:0] w1;    //: /sn:0 {0}(411,178)(#:330,178){1}
wire Cpy;    //: /sn:0 {0}(332,462)(332,452)(499,452)(499,-4){1}
wire [7:0] o3;    //: /sn:0 {0}(#:329,90)(427,90){1}
wire w17;    //: /sn:0 {0}(387,-4)(387,318){1}
wire w14;    //: /sn:0 {0}(435,85)(435,-4){1}
wire w11;    //: /sn:0 {0}(483,-4)(483,424)(352,424)(352,435){1}
wire w15;    //: /sn:0 {0}(419,-4)(419,173){1}
wire [7:0] o2;    //: /sn:0 {0}(#:322,383)(373,383){1}
wire w26;    //: /sn:0 {0}(403,250)(403,-4){1}
wire w9;    //: /sn:0 {0}(314,66)(314,67)(331,67)(331,57){1}
wire [7:0] o6;    //: /sn:0 {0}(379,323)(#:324,323){1}
//: enddecls

  _GGMUL8 #(124) g8 (.A(in2), .B(in1), .P(o5));   //: @(316,255) /sn:0 /R:1 /w:[ 11 13 0 ]
  _GGADD8 #(68, 70, 62, 64) g4 (.A(w6), .B(in1), .S(w1), .CI(w0), .CO(w4));   //: @(317,178) /sn:0 /R:1 /w:[ 0 9 1 0 0 ]
  _GGBUFIF8 #(4, 6) g47 (.Z(ALU_out), .I(in1), .E(Cpy));   //: @(330,467) /sn:0 /w:[ 33 29 0 ]
  //: GROUND g16 (w3) @(313,139) /sn:0 /w:[ 1 ]
  _GGADD8 #(68, 70, 62, 64) g3 (.A(in2), .B(in1), .S(o3), .CI(w9), .CO(w3));   //: @(316,90) /sn:0 /R:1 /w:[ 19 5 0 0 0 ]
  _GGBUFIF8 #(4, 6) g26 (.Z(ALU_out), .I(o3), .E(w14));   //: @(433,90) /sn:0 /w:[ 0 1 0 ]
  //: GROUND g17 (w4) @(345,223) /sn:0 /w:[ 1 ]
  //: LED g2 (w0) @(349,128) /sn:0 /w:[ 1 ] /type:0
  _GGBUFIF8 #(4, 6) g30 (.Z(ALU_out), .I(w37), .E(w18));   //: @(359,343) /sn:0 /w:[ 19 1 1 ]
  //: joint g23 (in1) @(131, 385) /w:[ 20 19 -1 22 ]
  //: joint g39 (ALU_out) @(650, 253) /w:[ -1 9 10 12 ]
  //: joint g24 (in1) @(131, 415) /w:[ 24 23 -1 26 ]
  //: IN g1 (in2) @(110,147) /sn:0 /w:[ 21 ]
  _GGBUFIF8 #(4, 6) g29 (.Z(ALU_out), .I(o6), .E(w17));   //: @(385,323) /sn:0 /w:[ 15 0 1 ]
  //: joint g18 (in1) @(131, 317) /w:[ 16 15 -1 18 ]
  dec4to16 g25 (.opc(opc), .o15(w23), .o14(w22), .o13(w21), .o12(w20), .o11(w19), .o10(w18), .o9(w17), .o8(w26), .o7(w15), .o6(w14), .o5(w13), .o4(w12), .o3(w11), .o2(Cpy), .o1(ST), .o0(LD));   //: @(275, -92) /sz:(272, 87) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 Bo1<0 Bo2<0 Bo3<0 Bo4<0 Bo5<0 Bo6<0 Bo7<1 Bo8<0 Bo9<1 Bo10<0 Bo11<0 Bo12<0 Bo13<1 Bo14<0 Bo15<0 ]
  //: joint g10 (in2) @(142, 194) /w:[ 14 -1 16 13 ]
  //: joint g49 (in1) @(122, 127) /w:[ 2 -1 1 28 ]
  //: joint g6 (in2) @(139, 147) /w:[ 18 -1 20 17 ]
  //: joint g35 (ALU_out) @(650, 411) /w:[ -1 25 26 28 ]
  //: joint g9 (in1) @(131, 162) /w:[ 8 7 -1 10 ]
  _GGNBUF8 #(2) g7 (.I(in2), .Z(w6));   //: @(192,194) /sn:0 /w:[ 15 1 ]
  _GGBUFIF8 #(4, 6) g31 (.Z(ALU_out), .I(o2), .E(w13));   //: @(379,383) /sn:0 /w:[ 23 1 1 ]
  //: joint g22 (in2) @(142, 380) /w:[ 2 4 -1 1 ]
  //: IN g45 (opc) @(532,-131) /sn:0 /R:3 /w:[ 1 ]
  //: joint g41 (ALU_out) @(651, 88) /w:[ -1 2 1 4 ]
  //: joint g36 (ALU_out) @(650, 381) /w:[ -1 21 22 24 ]
  _GGBUFIF8 #(4, 6) g33 (.Z(ALU_out), .I(o0), .E(w11));   //: @(350,440) /sn:0 /w:[ 31 1 1 ]
  //: OUT g42 (LD) @(547,42) /sn:0 /w:[ 1 ]
  //: joint g40 (ALU_out) @(650, 176) /w:[ -1 5 6 8 ]
  //: joint g12 (in1) @(131, 239) /w:[ 12 11 -1 14 ]
  //: OUT g34 (ALU_out) @(650,58) /sn:0 /R:1 /w:[ 3 ]
  _GGBUFIF8 #(4, 6) g28 (.Z(ALU_out), .I(o5), .E(w26));   //: @(401,255) /sn:0 /w:[ 11 1 0 ]
  //: joint g14 (in2) @(142, 349) /w:[ 6 8 -1 5 ]
  _GGDIV8 #(236, 236) g11 (.A(in2), .B(in1), .Q(o6), .R(w37));   //: @(311,333) /sn:0 /R:1 /w:[ 7 17 1 0 ]
  //: joint g5 (in1) @(131, 127) /w:[ 4 -1 3 6 ]
  _GGNBUF8 #(2) g21 (.I(in1), .Z(o0));   //: @(313,441) /sn:0 /w:[ 27 0 ]
  _GGAND2x8 #(6) g19 (.I0(in2), .I1(in1), .Z(o2));   //: @(312,383) /sn:0 /w:[ 3 21 0 ]
  _GGBUFIF8 #(4, 6) g32 (.Z(ALU_out), .I(o1), .E(w12));   //: @(362,413) /sn:0 /w:[ 27 1 1 ]
  _GGOR2x8 #(6) g20 (.I0(in2), .I1(in1), .Z(o1));   //: @(314,413) /sn:0 /w:[ 0 25 0 ]
  //: OUT g43 (ST) @(549,58) /sn:0 /w:[ 1 ]
  //: joint g38 (ALU_out) @(650, 321) /w:[ -1 13 14 16 ]
  //: LED g15 (w9) @(331,50) /sn:0 /w:[ 1 ] /type:0
  //: IN g0 (in1) @(109,127) /sn:0 /w:[ 0 ]
  //: joint g48 (ALU_out) @(650, 438) /w:[ -1 29 30 32 ]
  _GGBUFIF8 #(4, 6) g27 (.Z(ALU_out), .I(w1), .E(w15));   //: @(417,178) /sn:0 /w:[ 7 0 1 ]
  //: joint g37 (ALU_out) @(650, 341) /w:[ -1 17 18 20 ]
  //: joint g13 (in2) @(142, 271) /w:[ 10 12 -1 9 ]

endmodule
//: /netlistEnd

//: /netlistBegin Reg_file
module Reg_file(C, toRa, toRb, en_Rc, en_Ra, en_Rb, CLK, CLR, Ra_s, Rb_s, Rc_s);
//: interface  /sz:(124, 235) /bd:[ Ti0>C[7:0](61/124) Li0>CLR(190/235) Li1>CLK(172/235) Li2>Rb_s[1:0](121/235) Li3>en_Rb(105/235) Li4>Ra_s[1:0](54/235) Li5>en_Ra(28/235) Ri0>Rc_s[1:0](84/235) Ri1>en_Rc(112/235) Bo0<toRb[7:0](98/124) Bo1<toRa[7:0](21/124) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input en_Rc;    //: /sn:0 {0}(-49,-23)(-49,8)(-26,8){1}
input en_Rb;    //: /sn:0 {0}(498,-9)(498,29)(510,29){1}
input [1:0] Rc_s;    //: /sn:0 {0}(#:-2,-28)(-2,-5){1}
output [7:0] toRa;    //: /sn:0 {0}(#:397,301)(555,301)(555,251){1}
//: {2}(555,247)(555,231){3}
//: {4}(557,229)(#:581,229){5}
//: {6}(555,227)(555,195){7}
//: {8}(555,191)(555,135)(#:397,135){9}
//: {10}(553,193)(#:400,193){11}
//: {12}(553,249)(#:400,249){13}
input [1:0] Rb_s;    //: /sn:0 {0}(#:534,-6)(534,16){1}
input en_Ra;    //: /sn:0 {0}(406,-2)(406,33)(424,33){1}
input [1:0] Ra_s;    //: /sn:0 {0}(#:448,-1)(448,20){1}
input CLR;    //: /sn:0 {0}(311,45)(301,45)(301,58)(335,58)(335,109){1}
//: {2}(333,111)(320,111){3}
//: {4}(335,113)(335,171){5}
//: {6}(333,173)(324,173){7}
//: {8}(335,175)(335,226){9}
//: {10}(333,228)(326,228){11}
//: {12}(335,230)(335,275)(328,275){13}
input CLK;    //: /sn:0 {0}(88,278)(57,278)(57,233){1}
//: {2}(59,231)(63,231)(63,231)(88,231){3}
//: {4}(57,229)(57,177){5}
//: {6}(59,175)(77,175)(77,175)(88,175){7}
//: {8}(57,173)(57,115){9}
//: {10}(59,113)(77,113)(77,113)(88,113){11}
//: {12}(57,111)(57,56)(56,56)(56,7){13}
input [7:0] C;    //: /sn:0 {0}(#:150,5)(150,29){1}
//: {2}(152,31)(231,31)(#:231,106){3}
//: {4}(#:150,33)(150,152){5}
//: {6}(152,154)(232,154)(232,168){7}
//: {8}(150,156)(150,214){9}
//: {10}(152,216)(233,216)(233,224){11}
//: {12}(150,218)(150,258)(232,258)(232,271){13}
output [7:0] toRb;    //: /sn:0 {0}(#:500,420)(615,420)(615,394){1}
//: {2}(615,390)(615,375){3}
//: {4}(617,373)(#:635,373){5}
//: {6}(615,371)(615,360){7}
//: {8}(615,356)(615,330)(#:498,330){9}
//: {10}(613,358)(#:497,358){11}
//: {12}(613,392)(#:499,392){13}
supply0 w9;    //: /sn:0 {0}(271,286)(312,286){1}
//: {2}(314,284)(314,241){3}
//: {4}(314,237)(314,185){5}
//: {6}(314,181)(314,121)(270,121){7}
//: {8}(312,183)(271,183){9}
//: {10}(312,239)(272,239){11}
//: {12}(314,288)(314,328){13}
wire w16;    //: /sn:0 {0}(-20,24)(-20,283)(88,283){1}
wire w6;    //: /sn:0 {0}(16,24)(16,118)(88,118){1}
wire w13;    //: /sn:0 {0}(272,229)(294,229)(294,228)(310,228){1}
wire w7;    //: /sn:0 {0}(4,24)(4,180)(88,180){1}
wire w4;    //: /sn:0 {0}(109,116)(151,116)(151,116)(194,116){1}
wire w25;    //: /sn:0 {0}(528,45)(528,335)(489,335)(489,353){1}
wire w3;    //: /sn:0 {0}(270,111)(304,111){1}
wire [7:0] w0;    //: /sn:0 {0}(#:231,127)(231,135)(340,135){1}
//: {2}(344,135)(381,135){3}
//: {4}(#:342,137)(342,330)(482,330){5}
wire w22;    //: /sn:0 {0}(540,45)(540,369)(491,369)(491,387){1}
wire w20;    //: /sn:0 {0}(454,49)(454,229)(392,229)(392,244){1}
wire w29;    //: /sn:0 {0}(552,45)(552,400)(492,400)(492,415){1}
wire w19;    //: /sn:0 {0}(109,281)(155,281)(155,281)(195,281){1}
wire w18;    //: /sn:0 {0}(271,276)(290,276)(290,275)(312,275){1}
wire w12;    //: /sn:0 {0}(430,49)(430,115)(389,115)(389,130){1}
wire [7:0] w10;    //: /sn:0 {0}(#:233,245)(233,249)(354,249){1}
//: {2}(358,249)(384,249){3}
//: {4}(#:356,251)(356,392)(483,392){5}
wire w21;    //: /sn:0 {0}(466,49)(466,281)(389,281)(389,296){1}
wire w32;    //: /sn:0 {0}(516,45)(516,308)(490,308)(490,325){1}
wire w8;    //: /sn:0 {0}(271,173)(308,173){1}
wire w17;    //: /sn:0 {0}(442,49)(442,173)(392,173)(392,188){1}
wire w14;    //: /sn:0 {0}(109,234)(196,234){1}
wire w11;    //: /sn:0 {0}(-8,24)(-8,236)(88,236){1}
wire [7:0] w2;    //: /sn:0 {0}(#:232,189)(232,193)(346,193){1}
//: {2}(350,193)(384,193){3}
//: {4}(#:348,195)(348,358)(481,358){5}
wire [7:0] w15;    //: /sn:0 {0}(#:232,292)(232,301)(363,301){1}
//: {2}(367,301)(381,301){3}
//: {4}(#:365,303)(365,420)(484,420){5}
wire w26;    //: /sn:0 {0}(109,178)(156,178)(156,178)(195,178){1}
//: enddecls

  //: joint g8 (w9) @(314, 239) /w:[ -1 4 10 3 ]
  //: IN g4 (C) @(150,3) /sn:0 /R:3 /w:[ 0 ]
  //: joint g44 (C) @(150, 154) /w:[ 6 5 -1 8 ]
  _GGDECODER4 #(6, 6) g47 (.I(Rc_s), .E(en_Rc), .Z0(w6), .Z1(w7), .Z2(w11), .Z3(w16));   //: @(-2,8) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:1
  //: joint g16 (CLR) @(335, 228) /w:[ -1 9 10 12 ]
  _GGREG8 #(10, 10, 20) g3 (.Q(w15), .D(C), .EN(w9), .CLR(w18), .CK(w19));   //: @(232,281) /sn:0 /w:[ 0 13 0 0 1 ]
  //: OUT g17 (toRa) @(578,229) /sn:0 /w:[ 5 ]
  _GGBUFIF8 #(4, 6) g26 (.Z(toRa), .I(w15), .E(w21));   //: @(387,301) /sn:0 /w:[ 0 3 1 ]
  _GGREG8 #(10, 10, 20) g2 (.Q(w10), .D(C), .EN(w9), .CLR(w13), .CK(w14));   //: @(233,234) /sn:0 /w:[ 0 11 11 0 1 ]
  //: joint g23 (toRa) @(555, 193) /w:[ -1 8 10 7 ]
  _GGBUFIF8 #(4, 6) g30 (.Z(toRb), .I(w15), .E(w29));   //: @(490,420) /sn:0 /w:[ 0 5 1 ]
  _GGREG8 #(10, 10, 20) g1 (.Q(w2), .D(C), .EN(w9), .CLR(w8), .CK(w26));   //: @(232,178) /sn:0 /w:[ 0 7 9 0 1 ]
  _GGBUFIF8 #(4, 6) g24 (.Z(toRa), .I(w10), .E(w20));   //: @(390,249) /sn:0 /w:[ 13 3 1 ]
  //: joint g39 (toRb) @(615, 373) /w:[ 4 6 -1 3 ]
  _GGBUFIF8 #(4, 6) g29 (.Z(toRb), .I(w2), .E(w25));   //: @(487,358) /sn:0 /w:[ 11 5 1 ]
  //: joint g51 (CLK) @(57, 175) /w:[ 6 8 -1 5 ]
  //: OUT g18 (toRb) @(632,373) /sn:0 /w:[ 5 ]
  _GGNBUF #(2) g10 (.I(CLR), .Z(w18));   //: @(322,275) /sn:0 /R:2 /w:[ 13 1 ]
  //: joint g25 (toRa) @(555, 229) /w:[ 4 6 -1 3 ]
  _GGAND2 #(6) g49 (.I0(CLK), .I1(w7), .Z(w26));   //: @(99,178) /sn:0 /w:[ 7 1 0 ]
  //: joint g50 (CLK) @(57, 113) /w:[ 10 12 -1 9 ]
  //: GROUND g6 (w9) @(314,334) /sn:0 /w:[ 13 ]
  //: IN g56 (en_Rc) @(-49,-25) /sn:0 /R:3 /w:[ 0 ]
  //: joint g9 (w9) @(314, 183) /w:[ -1 6 8 5 ]
  //: joint g7 (w9) @(314, 286) /w:[ -1 2 1 12 ]
  //: joint g35 (w10) @(356, 249) /w:[ 2 -1 1 4 ]
  _GGBUFIF8 #(4, 6) g22 (.Z(toRa), .I(w2), .E(w17));   //: @(390,193) /sn:0 /w:[ 11 3 1 ]
  _GGBUFIF8 #(4, 6) g31 (.Z(toRb), .I(w0), .E(w32));   //: @(488,330) /sn:0 /w:[ 9 5 1 ]
  _GGAND2 #(6) g54 (.I0(CLK), .I1(w16), .Z(w19));   //: @(99,281) /sn:0 /w:[ 0 1 0 ]
  //: joint g33 (w2) @(348, 193) /w:[ 2 -1 1 4 ]
  //: joint g36 (w15) @(365, 301) /w:[ 2 -1 1 4 ]
  //: IN g41 (en_Ra) @(406,-4) /sn:0 /R:3 /w:[ 0 ]
  //: joint g45 (C) @(150, 216) /w:[ 10 9 -1 12 ]
  _GGAND2 #(6) g52 (.I0(CLK), .I1(w11), .Z(w14));   //: @(99,234) /sn:0 /w:[ 3 1 0 ]
  //: joint g40 (toRb) @(615, 392) /w:[ -1 2 12 1 ]
  //: IN g42 (en_Rb) @(498,-11) /sn:0 /R:3 /w:[ 0 ]
  _GGNBUF #(2) g12 (.I(CLR), .Z(w8));   //: @(318,173) /sn:0 /R:2 /w:[ 7 1 ]
  //: IN g46 (CLK) @(56,5) /sn:0 /R:3 /w:[ 13 ]
  _GGBUFIF8 #(4, 6) g28 (.Z(toRb), .I(w10), .E(w22));   //: @(489,392) /sn:0 /w:[ 13 5 1 ]
  _GGDECODER4 #(6, 6) g34 (.I(Ra_s), .E(en_Ra), .Z0(w12), .Z1(w17), .Z2(w20), .Z3(w21));   //: @(448,33) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  //: joint g14 (CLR) @(335, 111) /w:[ -1 1 2 4 ]
  _GGNBUF #(2) g11 (.I(CLR), .Z(w13));   //: @(320,228) /sn:0 /R:2 /w:[ 11 1 ]
  //: IN g5 (CLR) @(313,45) /sn:0 /R:2 /w:[ 0 ]
  //: IN g19 (Ra_s) @(448,-3) /sn:0 /R:3 /w:[ 0 ]
  _GGBUFIF8 #(4, 6) g21 (.Z(toRa), .I(w0), .E(w12));   //: @(387,135) /sn:0 /w:[ 9 3 1 ]
  //: IN g20 (Rb_s) @(534,-8) /sn:0 /R:3 /w:[ 0 ]
  //: joint g32 (w0) @(342, 135) /w:[ 2 -1 1 4 ]
  //: joint g15 (CLR) @(335, 173) /w:[ -1 5 6 8 ]
  _GGREG8 #(10, 10, 20) g0 (.Q(w0), .D(C), .EN(w9), .CLR(w3), .CK(w4));   //: @(231,116) /sn:0 /w:[ 0 3 7 0 1 ]
  //: joint g38 (toRb) @(615, 358) /w:[ -1 8 10 7 ]
  //: joint g43 (C) @(150, 31) /w:[ 2 1 -1 4 ]
  _GGAND2 #(6) g48 (.I0(CLK), .I1(w6), .Z(w4));   //: @(99,116) /sn:0 /w:[ 11 1 0 ]
  //: joint g27 (toRa) @(555, 249) /w:[ -1 2 12 1 ]
  _GGDECODER4 #(6, 6) g37 (.I(Rb_s), .E(en_Rb), .Z0(w32), .Z1(w25), .Z2(w22), .Z3(w29));   //: @(534,29) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  //: IN g55 (Rc_s) @(-2,-30) /sn:0 /R:3 /w:[ 0 ]
  //: joint g53 (CLK) @(57, 231) /w:[ 2 4 -1 1 ]
  _GGNBUF #(2) g13 (.I(CLR), .Z(w3));   //: @(314,111) /sn:0 /R:2 /w:[ 3 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin dec4to16
module dec4to16(o0, o8, o9, o15, o10, o2, o1, o14, o4, o6, o3, o13, o11, o12, o7, opc, o5);
//: interface  /sz:(87, 272) /bd:[ Li0>opc[3:0](16/272) Ro0<o0(16/272) Ro1<o1(32/272) Ro2<o2(48/272) Ro3<o3(64/272) Ro4<o4(80/272) Ro5<o5(96/272) Ro6<o6(112/272) Ro7<o7(128/272) Ro8<o8(144/272) Ro9<o9(160/272) Ro10<o10(176/272) Ro11<o11(192/272) Ro12<o12(208/272) Ro13<o13(224/272) Ro14<o14(240/272) Ro15<o15(256/272) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output o8;    //: /sn:0 {0}(527,105)(446,105)(446,107)(401,107){1}
output o1;    //: /sn:0 {0}(566,219)(479,219)(479,210)(400,210){1}
output o5;    //: /sn:0 {0}(563,181)(481,181)(481,183)(400,183){1}
output o10;    //: /sn:0 {0}(683,95)(673,95)(673,94)(401,94){1}
output o0;    //: /sn:0 {0}(519,235)(462,235)(462,217)(400,217){1}
input [3:0] opc;    //: /sn:0 {0}(#:159,259)(159,225){1}
//: {2}(159,224)(159,194){3}
//: {4}(159,193)(159,116){5}
//: {6}(159,115)(159,85){7}
//: {8}(159,84)(159,51){9}
output o9;    //: /sn:0 {0}(401,100)(489,100){1}
output o11;    //: /sn:0 {0}(712,87)(401,87){1}
output o7;    //: /sn:0 {0}(608,155)(462,155)(462,170)(400,170){1}
output o15;    //: /sn:0 {0}(659,61)(413,61)(413,60)(401,60){1}
output o12;    //: /sn:0 {0}(639,81)(407,81)(407,80)(401,80){1}
output o3;    //: /sn:0 {0}(547,197)(400,197){1}
output o4;    //: /sn:0 {0}(542,190)(400,190){1}
output o14;    //: /sn:0 {0}(617,67)(401,67){1}
output o13;    //: /sn:0 {0}(612,74)(401,74){1}
output o2;    //: /sn:0 {0}(400,203)(495,203)(495,209)(522,209){1}
output o6;    //: /sn:0 {0}(609,163)(525,163)(525,177)(400,177){1}
wire [2:0] w0;    //: /sn:0 {0}(163,85)(#:171,85)(171,84)(372,84){1}
wire [2:0] w10;    //: /sn:0 {0}(#:163,194)(371,194){1}
wire w21;    //: /sn:0 {0}(163,116)(267,116){1}
wire w1;    //: /sn:0 {0}(385,106)(385,116)(283,116){1}
wire w2;    //: /sn:0 {0}(163,225)(286,225){1}
wire w11;    //: /sn:0 {0}(302,225)(384,225)(384,216){1}
//: enddecls

  //: OUT g8 (o0) @(516,235) /sn:0 /w:[ 0 ]
  assign w21 = opc[3]; //: TAP g4 @(157,116) /sn:0 /R:2 /w:[ 0 5 6 ] /ss:1
  //: OUT g16 (o8) @(524,105) /sn:0 /w:[ 0 ]
  assign w0 = opc[2:0]; //: TAP g3 @(157,85) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:1
  //: OUT g17 (o9) @(486,100) /sn:0 /w:[ 1 ]
  _GGDECODER8 #(6, 6) g2 (.I(w10), .E(w11), .Z0(o0), .Z1(o1), .Z2(o2), .Z3(o3), .Z4(o4), .Z5(o5), .Z6(o6), .Z7(o7));   //: @(384,194) /sn:0 /R:1 /w:[ 1 1 1 1 0 1 1 1 1 1 ] /ss:0 /do:0
  //: OUT g23 (o15) @(656,61) /sn:0 /w:[ 0 ]
  _GGNBUF #(2) g24 (.I(w2), .Z(w11));   //: @(292,225) /sn:0 /w:[ 1 0 ]
  _GGDECODER8 #(6, 6) g1 (.I(w0), .E(w1), .Z0(o8), .Z1(o9), .Z2(o10), .Z3(o11), .Z4(o12), .Z5(o13), .Z6(o14), .Z7(o15));   //: @(385,84) /sn:0 /R:1 /w:[ 1 0 1 0 1 1 1 1 1 1 ] /ss:0 /do:0
  //: OUT g18 (o10) @(680,95) /sn:0 /w:[ 0 ]
  //: OUT g10 (o2) @(519,209) /sn:0 /w:[ 1 ]
  assign w10 = opc[2:0]; //: TAP g6 @(157,194) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  //: OUT g9 (o1) @(563,219) /sn:0 /w:[ 0 ]
  assign w2 = opc[3]; //: TAP g7 @(157,225) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: OUT g22 (o14) @(614,67) /sn:0 /w:[ 0 ]
  //: OUT g12 (o4) @(539,190) /sn:0 /w:[ 0 ]
  _GGBUF #(4) g5 (.I(w21), .Z(w1));   //: @(273,116) /sn:0 /w:[ 1 1 ]
  //: OUT g14 (o6) @(606,163) /sn:0 /w:[ 0 ]
  //: OUT g11 (o3) @(544,197) /sn:0 /w:[ 0 ]
  //: OUT g21 (o13) @(609,74) /sn:0 /w:[ 0 ]
  //: OUT g19 (o11) @(709,87) /sn:0 /w:[ 0 ]
  //: OUT g20 (o12) @(636,81) /sn:0 /w:[ 0 ]
  //: OUT g15 (o7) @(605,155) /sn:0 /w:[ 0 ]
  //: IN g0 (opc) @(159,261) /sn:0 /R:1 /w:[ 0 ]
  //: OUT g13 (o5) @(560,181) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

